`timescale 1ns / 1ps

/*
* This module is a uart receiver module. It receives the data coming from the external world
* and outputs the data.
*/
module uart_rx
#(
    parameter DATA_BITS = 8,    //Number of data bits to receieve via UART
              STOP_BITS = 1,    //Number of stop bits
              OVRSAMPLING = 16
)
(
    input logic clk, reset,
    input logic s_tick,                 //Input signal generated by the baudrate controller
    input logic rx,                     //Data coming into the UARt receiver
    output logic rx_done,               //Flag indicating reception is complete (all bits read)
    output logic [DATA_BITS-1:0] dout
);

/*********** Varibale declerations ***************/
localparam SB_TICKS = STOP_BITS * OVRSAMPLING;      //Number of ticks for the stop bits

//State Machine decleration
typedef enum {idle,                 //Initial starting state (when rx == 0 indicating start bit) switch states
              start,                //State to count the start bit ticks (7)
              data,                 //State to read the data
              stop} state_type;     //State to read the stop bits and signal completion

/*********** Signal Declerations ***************/
state_type state_reg, state_next;
logic [3:0] s_reg, s_next;                    //reg to keep track of smapling ticks (needs to count up to 15)
logic [2:0] n_reg, n_next;                    //reg to keep track of number of data bits recieved
logic [DATA_BITS-1:0] b_reg, b_next;          //reg to store the data coming into the receiever module

/********** UART Receiver Logic ****************/
always_ff @(posedge clk, posedge reset)
begin
    if(reset)
        begin
            state_reg <= idle;
            s_reg <= 0;
            n_reg <= 0;
            b_reg <= 0;
        end
    else
        begin
            state_reg <= state_next;
            s_reg <= s_next;
            n_reg <= n_next;
            b_reg <= b_next;
        end     
end

//Next State Logic
always_comb
begin
    //Default signals
    state_next = state_reg;
    s_next = s_reg;
    n_next = n_reg;
    b_next = b_reg;
    rx_done = 1'b0;
    //State Machine logic
    case(state_reg)
        idle:
        begin
            //If rx goes low (indicating start bit)
            if(~rx)
                begin
                    state_next = start;
                    s_next = 0;
                end        
        end
        start:
        begin
            //If tick from baud rate has been received 
            if(s_tick)
            begin
                //Once 7 tivks have been counted begin reading the data
                if(s_reg == 7)
                begin
                    state_next = data;
                    s_next = 0;
                    n_next = 0;
                end
                else
                    s_next = s_reg + 1;
            end                              
        end 
        data:
        begin
            if(s_tick)
            begin
                //if 15 ticks have been counted
                if(s_reg == 15)
                begin
                    s_next = 0;                         //Reset tick counter
                    b_next = {rx, b_reg[7:1]};          //Shift data into register
                    if(n_reg == (DATA_BITS - 1))        //If we have counted all the data bits
                        state_next = stop;
                    else
                        n_next = n_reg + 1;
                end
                else
                    s_next = s_reg + 1;
            end
        end 
        stop:
        begin
            if(s_tick)
            begin
                if(s_reg == (SB_TICKS-1))
                begin
                    state_next = idle;
                    rx_done = 1'b1;
                end
                else
                    s_next = s_reg + 1;
            end
        end     
    endcase
end

//Output logic
assign dout = b_reg;

endmodule
