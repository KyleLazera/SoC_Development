`timescale 1ns / 1ps

/*
* This module contains teh control logic for the spi slave that will interface with the SPi Master externally.
*/
module spi_slave
(
    input logic clk, reset,
    //Wrapper Interface
    output logic o_rx_done,                         //Flag indicating slave has complete a transaction
    output logic o_slave_rdy,                       //Flag indicating the slave is not undergoing a transaction
    output logic [7:0] o_mosi_byte,                 //The byte recieved by the Slave from the Master
    input logic [7:0] i_miso_byte,                  //This is the byte to transmit to the Master
    //SPI Interface Signals
    input logic i_spi_clk,                          //SPI Clock generated by SPI Master
    input logic i_spi_mosi,                         //MOSI generated by SPI Master
    input logic i_spi_cs_n,                         //Chip Select generated by SPI Master (active low)
    output logic o_spi_miso                         //MISO signal to ouput data to the SPI Master
);

//FSM States
typedef enum{idle,                  //Represents the initial phase before a transmission has begun
             mosi_sample,           //This phase is used to sample data on the rising edge
             miso_drive             //Used to transmit data on the falling edge
             }state_type;

/***** Signal Declarations ******/
state_type state_reg, state_next;
logic spi_clk_meta, spi_clk_reg, spi_clk;
logic spi_mosi_meta, spi_mosi_reg;
logic spi_cs_meta, spi_cs_reg;
logic r_edge_spi_clk, f_edge_spi_clk;
logic [2:0] bit_reg, bit_next;
logic [7:0] mosi_shift_reg, mosi_shift_next;
logic [7:0] miso_shift_reg, miso_shift_next;
logic rx_done;

/******** Synchronization Logic *********/
always_ff @(posedge clk) begin
    if(reset) begin
        spi_clk_meta <= 1'b0;
        spi_mosi_meta <= 1'b0;
        spi_cs_meta <= 1'b1;
        spi_clk_reg <= 1'b0;
        spi_mosi_reg <= 1'b0;
        spi_cs_reg <= 1'b1;
    end
    else begin
        spi_clk_meta <= i_spi_clk;
        spi_mosi_meta <= i_spi_mosi;
        spi_cs_meta <= i_spi_cs_n;
        spi_clk_reg <= spi_clk_meta;
        spi_mosi_reg <= spi_mosi_meta;
        spi_cs_reg <= spi_cs_meta;        
    end
end

/******** FSMD Logic for the Slave Reception/Sending **********/
//Synchrnonous Logic
always_ff @(posedge clk) begin
    if(reset) begin
        state_reg <= idle;
        spi_clk <= 1'b0;
        bit_reg <= 3'b111;
        mosi_shift_reg <= 8'b0;
        miso_shift_reg <= 8'b0;
    end
    else begin
        state_reg <= state_next;
        bit_reg <= bit_next;
        spi_clk <= spi_clk_reg;
        mosi_shift_reg <= mosi_shift_next;
        miso_shift_reg <= miso_shift_next;
    end
end

//Next-State Logic 
always_comb begin
    //Default Values - used to avoid inferred latches
    state_next = state_reg;
    bit_next = bit_reg;
    mosi_shift_next = mosi_shift_reg;
    miso_shift_next = miso_shift_reg;
    rx_done = 1'b0;
    o_slave_rdy = 1'b0;
    //FSM State Logic
    case(state_reg) 
        idle: begin
            o_slave_rdy = 1'b1;
            if(~spi_cs_reg) begin
                bit_next = 3'b111;
                o_slave_rdy = 1'b0;
                mosi_shift_next = 8'b0;
                miso_shift_next = i_miso_byte;
                state_next = mosi_sample;
            end
        end        
        mosi_sample : begin
            //If cs is low and rising edge of spi slock is detected
            if(r_edge_spi_clk && ~spi_cs_reg) begin
                //shift the MOSI signal into the mosi shift reg
                mosi_shift_next = {mosi_shift_reg, spi_mosi_reg};
                state_next = miso_drive;
            end
        end        
        miso_drive : begin
            //If there is a falling edge and chip select is active
            if(f_edge_spi_clk && ~spi_cs_reg) begin
                //Shift the mosi shift reg to the left by 1 so the MSB can be output
                miso_shift_next = {miso_shift_reg[6:0], 1'b0};
                if(bit_reg == 3'b0) begin
                    bit_next = 3'b111;
                    rx_done = 1'b1;
                    state_next = idle;
                end
                else begin
                    bit_next = bit_reg - 1;
                    state_next = mosi_sample;
                end           
            end
        end
    endcase
end

//Rising & Falling edge detection Signals
assign r_edge_spi_clk = ~spi_clk & spi_clk_reg;
assign f_edge_spi_clk = spi_clk & ~spi_clk_reg;

//Output Logic
assign o_rx_done = rx_done;
assign o_mosi_byte = mosi_shift_reg;
assign o_spi_miso = miso_shift_reg[7];

endmodule
