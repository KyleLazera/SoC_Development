`timescale 1ns / 1ps


/* This module is used to test the PWM module using a large variety of possible values on one of the output channels. It is a self-checking testbench that
* utilizes OOP principles. The architecutre of the Testbench is as follows:
* pwm_driver : This class drives generated values to the actual hardware design via a virtual interface
* pwm_monitor : This class monitors the hardware via teh virtual interface and does some basic calculations to determine what the
                diviosr and duty cycle are based purley on the output of the hardware
* scoreboard : This class compares teh calculated values from the monitor to the expected values which are generated by the driver.
                This class also outputs the final scoreboard letting the suer know if all transmissions were succesful
* environemnt : This class encapsulates the driver, monitor and scoreboard into a singular environemnt that can be reused
* test : This class is used to generate the signals that are sent to the driver. This class encapsulates the environment and interfaces with the
        top level testbench.
*/
module pwm_tb_top;

    logic clk, reset;
    //Inst clock with 10 ns period
    always #5 clk = ~clk;
    //Init the virtual interface
    pwm_if  pwm_vif(clk, reset);
    
    //Module inst
    pwm_core #(.OUT_PORTS(6), .RES(8)) pwm_dut(.clk(clk), .reset(reset), .cs(pwm_vif.cs), .read(pwm_vif.read), .write(pwm_vif.write),
                                               .reg_addr(pwm_vif.reg_addr), .wr_data(pwm_vif.wr_data), .rd_data(pwm_vif.rd_data), 
                                               .pwm_out(pwm_vif.pwm_out));
                                               
    //Test Instance
    pwm_test default_test;
    
    initial begin
        clk = 0;
        
        //Reset the circuit
        reset = 1'b1;
        #10;
        reset = 1'b0;
        
        default_test = new(pwm_vif);
        default_test.env.vif = pwm_vif;
        default_test.main();
        
        #200;
        $finish;
    end


endmodule
